// ============================================================================
// File: hazard_unit.v
// Description: Hazard Detection Unit for ARM Cortex-A9 Pipeline
// Course: 05_ARM_Cortex_A9 - AI4ICLearning
// ============================================================================

`include "defines.vh"

module hazard_unit (
    // ========================================================================
    // 时钟与复位
    // ========================================================================
    input  wire                     clk,
    input  wire                     rst_n,
    
    // ========================================================================
    // ID 阶段信息
    // ========================================================================
    input  wire [3:0]               id_rn,          // 源寄存器 1
    input  wire [3:0]               id_rm,          // 源寄存器 2
    input  wire [3:0]               id_rs,          // 移位寄存器
    input  wire                     id_branch,      // 分支指令
    
    // ========================================================================
    // EX 阶段信息
    // ========================================================================
    input  wire [3:0]               ex_rd,          // 目的寄存器
    input  wire                     ex_mem_read,    // Load 指令
    input  wire                     ex_reg_write,   // 寄存器写使能
    
    // ========================================================================
    // MEM 阶段信息
    // ========================================================================
    input  wire [3:0]               mem_rd,         // 目的寄存器
    input  wire                     mem_reg_write,  // 寄存器写使能
    
    // ========================================================================
    // 分支信号
    // ========================================================================
    input  wire                     branch_taken,   // 分支被执行
    
    // ========================================================================
    // 控制输出
    // ========================================================================
    output reg                      stall_if,       // IF 阶段暂停
    output reg                      stall_id,       // ID 阶段暂停
    output reg                      flush_if,       // IF 阶段冲刷
    output reg                      flush_id,       // ID 阶段冲刷
    output reg                      flush_ex        // EX 阶段冲刷
);

    // ========================================================================
    // Load-Use 冒险检测
    // ========================================================================
    
    // 检测 EX 阶段的 Load 指令是否与 ID 阶段指令存在依赖
    wire load_use_hazard;
    
    assign load_use_hazard = ex_mem_read && ex_reg_write && (ex_rd != 4'd0) &&
                             ((ex_rd == id_rn) || (ex_rd == id_rm) || (ex_rd == id_rs));
    
    // ========================================================================
    // 分支冒险检测
    // ========================================================================
    
    // 分支目标在 EX 阶段确定，需要冲刷 IF 和 ID 阶段
    wire branch_hazard;
    
    assign branch_hazard = branch_taken;
    
    // ========================================================================
    // 控制信号生成
    // ========================================================================
    
    always @(*) begin
        // 默认值：不暂停，不冲刷
        stall_if = 1'b0;
        stall_id = 1'b0;
        flush_if = 1'b0;
        flush_id = 1'b0;
        flush_ex = 1'b0;
        
        // --------------------------------------------------------------------
        // Load-Use 冒险处理
        // 暂停 IF 和 ID，在 EX 插入气泡
        // --------------------------------------------------------------------
        if (load_use_hazard) begin
            stall_if = 1'b1;
            stall_id = 1'b1;
            flush_ex = 1'b1;  // 插入 NOP
        end
        
        // --------------------------------------------------------------------
        // 分支冒险处理
        // 冲刷 IF 和 ID 阶段（分支已在 EX 阶段确定）
        // --------------------------------------------------------------------
        if (branch_hazard) begin
            flush_if = 1'b1;
            flush_id = 1'b1;
            // 如果同时存在 Load-Use 冒险，分支优先
            stall_if = 1'b0;
            stall_id = 1'b0;
        end
    end

endmodule
