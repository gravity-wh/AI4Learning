// ============================================================================
// File: forwarding_unit.v
// Description: Data Forwarding Unit for ARM Cortex-A9 Pipeline
// Course: 05_ARM_Cortex_A9 - AI4ICLearning
// ============================================================================

`include "defines.vh"

module forwarding_unit (
    // ========================================================================
    // EX 阶段源寄存器
    // ========================================================================
    input  wire [3:0]               ex_rn,          // Operand A 源寄存器
    input  wire [3:0]               ex_rm,          // Operand B 源寄存器
    
    // ========================================================================
    // MEM 阶段信息
    // ========================================================================
    input  wire [3:0]               mem_rd,         // MEM 目的寄存器
    input  wire                     mem_reg_write,  // MEM 寄存器写使能
    
    // ========================================================================
    // WB 阶段信息
    // ========================================================================
    input  wire [3:0]               wb_rd,          // WB 目的寄存器
    input  wire                     wb_reg_write,   // WB 寄存器写使能
    
    // ========================================================================
    // 前递控制输出
    // ========================================================================
    output reg  [1:0]               forward_a,      // Operand A 前递选择
    output reg  [1:0]               forward_b       // Operand B 前递选择
);

    // ========================================================================
    // 前递逻辑 - Operand A (Rn)
    // ========================================================================
    
    always @(*) begin
        // 默认不前递，使用寄存器文件数据
        forward_a = `FWD_NONE;
        
        // MEM 冒险检测 (MEM→EX 前递，优先级更高)
        // 条件：MEM 阶段写入的寄存器正是 EX 阶段需要的源寄存器
        if (mem_reg_write && 
            (mem_rd != 4'd0) &&     // R0 不需要前递（假设 R0 恒为 0）
            (mem_rd != 4'd15) &&    // PC 特殊处理
            (mem_rd == ex_rn)) begin
            forward_a = `FWD_MEM;
        end
        // WB 冒险检测 (WB→EX 前递)
        // 条件：WB 阶段写入的寄存器正是 EX 阶段需要的源寄存器
        //       且 MEM 阶段没有写同一个寄存器
        else if (wb_reg_write && 
                 (wb_rd != 4'd0) &&
                 (wb_rd != 4'd15) &&
                 (wb_rd == ex_rn)) begin
            forward_a = `FWD_WB;
        end
    end
    
    // ========================================================================
    // 前递逻辑 - Operand B (Rm)
    // ========================================================================
    
    always @(*) begin
        // 默认不前递
        forward_b = `FWD_NONE;
        
        // MEM 冒险检测
        if (mem_reg_write && 
            (mem_rd != 4'd0) &&
            (mem_rd != 4'd15) &&
            (mem_rd == ex_rm)) begin
            forward_b = `FWD_MEM;
        end
        // WB 冒险检测
        else if (wb_reg_write && 
                 (wb_rd != 4'd0) &&
                 (wb_rd != 4'd15) &&
                 (wb_rd == ex_rm)) begin
            forward_b = `FWD_WB;
        end
    end

endmodule
